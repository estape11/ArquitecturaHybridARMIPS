module Test(input logic [31:0] in, output logic [2:0] out);
	assign out=in[25:23];
endmodule 